pll108MHz_inst : pll108MHz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
